module Alu (data1, data2, select, result);
  input[7:0] data1, data2;
  input[2:0] select;
  output [7:0] result;

  //TODO: Instantiate sub-units 
  
endmodule