module Task1;
endmodule




